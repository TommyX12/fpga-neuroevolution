
module main();
    
endmodule
