module draw_background(
	input start,
	input clock,
	output drawing,
	output x,
	output y,
	output colour,	// WE'RE CANADIAN
	output plot
	);
	
	
	
	always @(posedge clock) begin
		
	end

endmodule
